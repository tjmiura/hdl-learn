/* AND2 */

module AND2 ( A, B, X );

input A, B;
output X;

  and AAA (X, A, B);

endmodule
